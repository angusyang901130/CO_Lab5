`timescale 1ns/1ps
module Pipeline_CPU(
    clk_i,
    rst_i
);

//I/O port
input         clk_i;
input         rst_i;

//Internal Signals
wire [31:0] PC_i; // input in IF, output in IF
wire [31:0] PC_o; // input in IF, output in IF, input in IF/ID
wire [31:0] MUXMemtoReg_o;
wire [31:0] ALUResult;
wire [31:0] MUXALUSrc_o;
wire [31:0] Decoder_o;
wire [31:0] RSdata_o;
wire [31:0] RTdata_o;
wire [31:0] Imm_Gen_o;
wire [31:0] ALUSrc1_o;
wire [31:0] ALUSrc2_o;
wire [7:0]  MUX_control_o;

wire [31:0] PC_Add_Immediate; // input in IF
wire [1:0] ALUOp;
wire PC_write; // input in IF
wire ALUSrc;
wire RegWrite;
wire Branch;
wire MUXControl; // generated by hazard detection unit
wire Jump;
wire [31:0] SL1_o;
wire [3:0] ALU_Ctrl_o;
wire ALU_zero;
wire Branch_zero;
wire MUXPCSrc; // input in IF
wire [31:0] DM_o;
wire MemtoReg, MemRead, MemWrite;
wire [1:0] ForwardA;    // output in EXE
wire [1:0] ForwardB;    // output in EXE
wire [31:0] PC_Add4;  // input in IF


//Pipeline Register Signals
//IFID
wire [31:0] IFID_PC_o;
wire [31:0] IFID_Instr_o;
wire IFID_Write;
wire IFID_Flush; 
wire [31:0]IFID_PC_Add4_o;

//IDEXE
wire [31:0] IDEXE_Instr_o;
wire [2:0] IDEXE_WB_o;
wire [1:0] IDEXE_Mem_o;
wire [2:0] IDEXE_Exe_o;
wire [31:0] IDEXE_PC_o;
wire [31:0] IDEXE_RSdata_o;
wire [31:0] IDEXE_RTdata_o;
wire [31:0] IDEXE_ImmGen_o;
wire [3:0] IDEXE_Instr_30_14_12_o;
wire [4:0] IDEXE_Instr_11_7_o;
wire [31:0]IDEXE_PC_add4_o;

//EXEMEM
wire [31:0] EXEMEM_Instr_o;
wire [2:0] EXEMEM_WB_o;
wire [1:0] EXEMEM_Mem_o;
wire [31:0] EXEMEM_PCsum_o;
wire EXEMEM_Zero_o;
wire [31:0] EXEMEM_ALUResult_o;
wire [31:0] EXEMEM_RTdata_o;
wire [4:0]  EXEMEM_Instr_11_7_o;
wire [31:0] EXEMEM_PC_Add4_o;

//MEMWB
wire [2:0] MEMWB_WB_o;
wire [31:0] MEMWB_DM_o;
wire [31:0] MEMWB_ALUresult_o;
wire [4:0]  MEMWB_Instr_11_7_o;
wire [31:0] MEMWB_PC_Add4_o;

// wire
wire [31:0] imm_4 = 4; // input in IF
wire [31:0] instr; // output in IF, input 

// IF 
MUX_2to1 MUX_PCSrc(
    .data0_i(PC_Add4),
    .data1_i(PC_Add_Immediate),
    .select_i(MUXPCSrc),
    .data_o(PC_i)
);

ProgramCounter PC(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .PCwrite(PC_write),
    .pc_i(PC_i),
    .pc_o(PC_o)
);

Adder PC_plus_4_Adder(
    .src1_i(PC_o),
    .src2_i(imm_4),
    .sum_o(PC_Add4)
);

Instr_Memory IM(
    .addr_i(PC_o),
    .instr_o(instr)
);

IFID_register IFtoID(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .flush(IFID_Flush),
    .IFID_write(IFID_Write),
    .address_i(PC_o),
    .instr_i(instr),
    .pc_add4_i(PC_Add4),
    .address_o(IFID_PC_o),
    .instr_o(IFID_Instr_o),
    .pc_add4_o(IFID_PC_Add4_o)
);

// ID
Hazard_detection Hazard_detection_obj(

);

MUX_2to1 MUX_control(
    
);

Decoder Decoder(
);

Reg_File RF(
);

Imm_Gen ImmGen(
);

Shift_Left_1 SL1(
);

Adder Branch_Adder(
);

IDEXE_register IDtoEXE(
);

// EXE
MUX_2to1 MUX_ALUSrc(
    .data0_i(),
    .data1_i(),
    .select_i(),
    .data_o()
);

ForwardingUnit FWUnit(
    .IDEXE_RS1(),
    .IDEXE_RS2(),
    .EXEMEM_RD(),
    .MEMWB_RD(),
    .EXEMEM_RegWrite(),
    .MEMWB_RegWrite(),
    .ForwardA(ForwardA),
    .ForwardB(ForwardB)
);

MUX_3to1 MUX_ALU_src1(
    .data0_i(),
    .data1_i(),
    .data2_i(),
    .select_i(ForwardA),
    .data_o()
);

MUX_3to1 MUX_ALU_src2(
    .data0_i(),
    .data1_i(),
    .data2_i(),
    .select_i(ForwardB),
    .data_o()
);

ALU_Ctrl ALU_Ctrl(
    .instr(),
    .ALUOp(),
    .ALU_Ctrl_o()
);

alu alu(
    .rst_n(rst_i),
    .src1(),
    .src2(),
    .ALU_control(),
    .result(),
    .Zero()
);

EXEMEM_register EXEtoMEM(
    .clk_i(clk_i),
	.rst_i(),
	.instr_i(),
	.WB_i(),
	.Mem_i(),
	.zero_i(),
	.alu_ans_i(),
	.rtdata_i(),
	.WBreg_i(),
	.pc_add4_i(),
	.instr_o(),
	.WB_o(),
	.Mem_o(),
	.zero_o(),
	.alu_ans_o(),
	.rtdata_o(),
	.WBreg_o(),
	.pc_add4_o()
);

// MEM
Data_Memory Data_Memory(
    .clk_i(clk_i),
    .addr_i(),
    .data_i(),
    .MemRead_i(),
    .MemWrite_i(),
    .data_o()
);

MEMWB_register MEMtoWB(
    .clk_i(clk_i),
    .rst_i(),
    .WB_i(),
    .DM_i(),
    .alu_ans_i(),
    .WBreg_i(),
    .pc_add4_i(),
    .WB_o(),
    .DM_o(),
    .alu_ans_o(),
    .WBreg_o(),
    .pc_add4_o()
);

// WB
MUX_3to1 MUX_MemtoReg(
    .data0_i(),
    .data1_i(),
    .data2_i(),
    .select_i(),
    .data_o()
);

endmodule



